// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CLK_ST_CHKR_SV__
`define __UVME_CLK_ST_CHKR_SV__


/**
 * TODO Describe uvme_clk_st_chkr
 */
module uvme_clk_st_chkr (
      uvma_clk_if  active_if,
      uvma_clk_if  passive_if
);
   
   // TODO Add assertions to uvme_clk_st_chkr
   
endmodule : uvme_clk_st_chkr


`endif // __UVME_CLK_ST_CHKR_SV__
