// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CLK_IF_CHKR_SV__
`define __UVMA_CLK_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_clk_if.
 */
module uvma_clk_if_chkr(
   uvma_clk_if  clk_if
);
   
   // TODO Add assertions to uvma_clk_if_chkr
   
endmodule : uvma_clk_if_chkr


`endif // __UVMA_CLK_IF_CHKR_SV__
