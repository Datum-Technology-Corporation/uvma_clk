// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CLK_ST_DUT_CHKR_SV__
`define __UVMT_CLK_ST_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for Clock VIP
 * Self-Testing DUT wrapper (uvmt_clk_st_dut_wrap).
 */
module uvmt_clk_st_dut_chkr(
   uvma_clk_if  active_if,
   uvma_clk_if  passive_if
);
   
   // TODO Add assertions to uvmt_clk_st_dut_chkr
   
endmodule : uvmt_clk_st_dut_chkr


`endif // __UVMT_CLK_ST_DUT_CHKR_SV__
