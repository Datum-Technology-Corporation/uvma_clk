// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CLK_ST_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_CLK_ST_BASE_TEST_WORKAROUNDS_SV__


// This file should be empty by the end of the project


`endif // __UVMT_CLK_ST_BASE_TEST_WORKAROUNDS_SV__
