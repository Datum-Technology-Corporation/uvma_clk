// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CLK_MACROS_SV__
`define __UVMA_CLK_MACROS_SV__


`define UVMA_CLK_DEFAULT_FREQUENCY   100_000_000
`define UVMA_CLK_DEFAULT_DUTY_CYCLE           50


`endif // __UVMA_CLK_MACROS_SV__
